magic
tech sky130A
magscale 1 2
timestamp 1624040041
<< obsli1 >>
rect 1104 85 238832 197489
<< obsm1 >>
rect 290 8 239738 197520
<< metal2 >>
rect 1030 199200 1086 200000
rect 3054 199200 3110 200000
rect 5170 199200 5226 200000
rect 7286 199200 7342 200000
rect 9310 199200 9366 200000
rect 11426 199200 11482 200000
rect 13542 199200 13598 200000
rect 15566 199200 15622 200000
rect 17682 199200 17738 200000
rect 19798 199200 19854 200000
rect 21822 199200 21878 200000
rect 23938 199200 23994 200000
rect 26054 199200 26110 200000
rect 28078 199200 28134 200000
rect 30194 199200 30250 200000
rect 32310 199200 32366 200000
rect 34334 199200 34390 200000
rect 36450 199200 36506 200000
rect 38566 199200 38622 200000
rect 40682 199200 40738 200000
rect 42706 199200 42762 200000
rect 44822 199200 44878 200000
rect 46938 199200 46994 200000
rect 48962 199200 49018 200000
rect 51078 199200 51134 200000
rect 53194 199200 53250 200000
rect 55218 199200 55274 200000
rect 57334 199200 57390 200000
rect 59450 199200 59506 200000
rect 61474 199200 61530 200000
rect 63590 199200 63646 200000
rect 65706 199200 65762 200000
rect 67730 199200 67786 200000
rect 69846 199200 69902 200000
rect 71962 199200 72018 200000
rect 74078 199200 74134 200000
rect 76102 199200 76158 200000
rect 78218 199200 78274 200000
rect 80334 199200 80390 200000
rect 82358 199200 82414 200000
rect 84474 199200 84530 200000
rect 86590 199200 86646 200000
rect 88614 199200 88670 200000
rect 90730 199200 90786 200000
rect 92846 199200 92902 200000
rect 94870 199200 94926 200000
rect 96986 199200 97042 200000
rect 99102 199200 99158 200000
rect 101126 199200 101182 200000
rect 103242 199200 103298 200000
rect 105358 199200 105414 200000
rect 107474 199200 107530 200000
rect 109498 199200 109554 200000
rect 111614 199200 111670 200000
rect 113730 199200 113786 200000
rect 115754 199200 115810 200000
rect 117870 199200 117926 200000
rect 119986 199200 120042 200000
rect 122010 199200 122066 200000
rect 124126 199200 124182 200000
rect 126242 199200 126298 200000
rect 128266 199200 128322 200000
rect 130382 199200 130438 200000
rect 132498 199200 132554 200000
rect 134522 199200 134578 200000
rect 136638 199200 136694 200000
rect 138754 199200 138810 200000
rect 140870 199200 140926 200000
rect 142894 199200 142950 200000
rect 145010 199200 145066 200000
rect 147126 199200 147182 200000
rect 149150 199200 149206 200000
rect 151266 199200 151322 200000
rect 153382 199200 153438 200000
rect 155406 199200 155462 200000
rect 157522 199200 157578 200000
rect 159638 199200 159694 200000
rect 161662 199200 161718 200000
rect 163778 199200 163834 200000
rect 165894 199200 165950 200000
rect 167918 199200 167974 200000
rect 170034 199200 170090 200000
rect 172150 199200 172206 200000
rect 174266 199200 174322 200000
rect 176290 199200 176346 200000
rect 178406 199200 178462 200000
rect 180522 199200 180578 200000
rect 182546 199200 182602 200000
rect 184662 199200 184718 200000
rect 186778 199200 186834 200000
rect 188802 199200 188858 200000
rect 190918 199200 190974 200000
rect 193034 199200 193090 200000
rect 195058 199200 195114 200000
rect 197174 199200 197230 200000
rect 199290 199200 199346 200000
rect 201314 199200 201370 200000
rect 203430 199200 203486 200000
rect 205546 199200 205602 200000
rect 207662 199200 207718 200000
rect 209686 199200 209742 200000
rect 211802 199200 211858 200000
rect 213918 199200 213974 200000
rect 215942 199200 215998 200000
rect 218058 199200 218114 200000
rect 220174 199200 220230 200000
rect 222198 199200 222254 200000
rect 224314 199200 224370 200000
rect 226430 199200 226486 200000
rect 228454 199200 228510 200000
rect 230570 199200 230626 200000
rect 232686 199200 232742 200000
rect 234710 199200 234766 200000
rect 236826 199200 236882 200000
rect 238942 199200 238998 200000
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2134 0 2190 800
rect 2594 0 2650 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6550 0 6606 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 8022 0 8078 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9954 0 10010 800
rect 10414 0 10470 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12898 0 12954 800
rect 13358 0 13414 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15842 0 15898 800
rect 16302 0 16358 800
rect 16762 0 16818 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18694 0 18750 800
rect 19246 0 19302 800
rect 19706 0 19762 800
rect 20166 0 20222 800
rect 20718 0 20774 800
rect 21178 0 21234 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22650 0 22706 800
rect 23110 0 23166 800
rect 23662 0 23718 800
rect 24122 0 24178 800
rect 24582 0 24638 800
rect 25042 0 25098 800
rect 25594 0 25650 800
rect 26054 0 26110 800
rect 26514 0 26570 800
rect 27066 0 27122 800
rect 27526 0 27582 800
rect 27986 0 28042 800
rect 28538 0 28594 800
rect 28998 0 29054 800
rect 29458 0 29514 800
rect 30010 0 30066 800
rect 30470 0 30526 800
rect 30930 0 30986 800
rect 31482 0 31538 800
rect 31942 0 31998 800
rect 32402 0 32458 800
rect 32954 0 33010 800
rect 33414 0 33470 800
rect 33874 0 33930 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35346 0 35402 800
rect 35806 0 35862 800
rect 36358 0 36414 800
rect 36818 0 36874 800
rect 37278 0 37334 800
rect 37830 0 37886 800
rect 38290 0 38346 800
rect 38750 0 38806 800
rect 39302 0 39358 800
rect 39762 0 39818 800
rect 40222 0 40278 800
rect 40774 0 40830 800
rect 41234 0 41290 800
rect 41694 0 41750 800
rect 42154 0 42210 800
rect 42706 0 42762 800
rect 43166 0 43222 800
rect 43626 0 43682 800
rect 44178 0 44234 800
rect 44638 0 44694 800
rect 45098 0 45154 800
rect 45650 0 45706 800
rect 46110 0 46166 800
rect 46570 0 46626 800
rect 47122 0 47178 800
rect 47582 0 47638 800
rect 48042 0 48098 800
rect 48594 0 48650 800
rect 49054 0 49110 800
rect 49514 0 49570 800
rect 49974 0 50030 800
rect 50526 0 50582 800
rect 50986 0 51042 800
rect 51446 0 51502 800
rect 51998 0 52054 800
rect 52458 0 52514 800
rect 52918 0 52974 800
rect 53470 0 53526 800
rect 53930 0 53986 800
rect 54390 0 54446 800
rect 54942 0 54998 800
rect 55402 0 55458 800
rect 55862 0 55918 800
rect 56414 0 56470 800
rect 56874 0 56930 800
rect 57334 0 57390 800
rect 57886 0 57942 800
rect 58346 0 58402 800
rect 58806 0 58862 800
rect 59266 0 59322 800
rect 59818 0 59874 800
rect 60278 0 60334 800
rect 60738 0 60794 800
rect 61290 0 61346 800
rect 61750 0 61806 800
rect 62210 0 62266 800
rect 62762 0 62818 800
rect 63222 0 63278 800
rect 63682 0 63738 800
rect 64234 0 64290 800
rect 64694 0 64750 800
rect 65154 0 65210 800
rect 65706 0 65762 800
rect 66166 0 66222 800
rect 66626 0 66682 800
rect 67086 0 67142 800
rect 67638 0 67694 800
rect 68098 0 68154 800
rect 68558 0 68614 800
rect 69110 0 69166 800
rect 69570 0 69626 800
rect 70030 0 70086 800
rect 70582 0 70638 800
rect 71042 0 71098 800
rect 71502 0 71558 800
rect 72054 0 72110 800
rect 72514 0 72570 800
rect 72974 0 73030 800
rect 73526 0 73582 800
rect 73986 0 74042 800
rect 74446 0 74502 800
rect 74906 0 74962 800
rect 75458 0 75514 800
rect 75918 0 75974 800
rect 76378 0 76434 800
rect 76930 0 76986 800
rect 77390 0 77446 800
rect 77850 0 77906 800
rect 78402 0 78458 800
rect 78862 0 78918 800
rect 79322 0 79378 800
rect 79874 0 79930 800
rect 80334 0 80390 800
rect 80794 0 80850 800
rect 81346 0 81402 800
rect 81806 0 81862 800
rect 82266 0 82322 800
rect 82818 0 82874 800
rect 83278 0 83334 800
rect 83738 0 83794 800
rect 84198 0 84254 800
rect 84750 0 84806 800
rect 85210 0 85266 800
rect 85670 0 85726 800
rect 86222 0 86278 800
rect 86682 0 86738 800
rect 87142 0 87198 800
rect 87694 0 87750 800
rect 88154 0 88210 800
rect 88614 0 88670 800
rect 89166 0 89222 800
rect 89626 0 89682 800
rect 90086 0 90142 800
rect 90638 0 90694 800
rect 91098 0 91154 800
rect 91558 0 91614 800
rect 92018 0 92074 800
rect 92570 0 92626 800
rect 93030 0 93086 800
rect 93490 0 93546 800
rect 94042 0 94098 800
rect 94502 0 94558 800
rect 94962 0 95018 800
rect 95514 0 95570 800
rect 95974 0 96030 800
rect 96434 0 96490 800
rect 96986 0 97042 800
rect 97446 0 97502 800
rect 97906 0 97962 800
rect 98458 0 98514 800
rect 98918 0 98974 800
rect 99378 0 99434 800
rect 99838 0 99894 800
rect 100390 0 100446 800
rect 100850 0 100906 800
rect 101310 0 101366 800
rect 101862 0 101918 800
rect 102322 0 102378 800
rect 102782 0 102838 800
rect 103334 0 103390 800
rect 103794 0 103850 800
rect 104254 0 104310 800
rect 104806 0 104862 800
rect 105266 0 105322 800
rect 105726 0 105782 800
rect 106278 0 106334 800
rect 106738 0 106794 800
rect 107198 0 107254 800
rect 107750 0 107806 800
rect 108210 0 108266 800
rect 108670 0 108726 800
rect 109130 0 109186 800
rect 109682 0 109738 800
rect 110142 0 110198 800
rect 110602 0 110658 800
rect 111154 0 111210 800
rect 111614 0 111670 800
rect 112074 0 112130 800
rect 112626 0 112682 800
rect 113086 0 113142 800
rect 113546 0 113602 800
rect 114098 0 114154 800
rect 114558 0 114614 800
rect 115018 0 115074 800
rect 115570 0 115626 800
rect 116030 0 116086 800
rect 116490 0 116546 800
rect 116950 0 117006 800
rect 117502 0 117558 800
rect 117962 0 118018 800
rect 118422 0 118478 800
rect 118974 0 119030 800
rect 119434 0 119490 800
rect 119894 0 119950 800
rect 120446 0 120502 800
rect 120906 0 120962 800
rect 121366 0 121422 800
rect 121918 0 121974 800
rect 122378 0 122434 800
rect 122838 0 122894 800
rect 123390 0 123446 800
rect 123850 0 123906 800
rect 124310 0 124366 800
rect 124770 0 124826 800
rect 125322 0 125378 800
rect 125782 0 125838 800
rect 126242 0 126298 800
rect 126794 0 126850 800
rect 127254 0 127310 800
rect 127714 0 127770 800
rect 128266 0 128322 800
rect 128726 0 128782 800
rect 129186 0 129242 800
rect 129738 0 129794 800
rect 130198 0 130254 800
rect 130658 0 130714 800
rect 131210 0 131266 800
rect 131670 0 131726 800
rect 132130 0 132186 800
rect 132590 0 132646 800
rect 133142 0 133198 800
rect 133602 0 133658 800
rect 134062 0 134118 800
rect 134614 0 134670 800
rect 135074 0 135130 800
rect 135534 0 135590 800
rect 136086 0 136142 800
rect 136546 0 136602 800
rect 137006 0 137062 800
rect 137558 0 137614 800
rect 138018 0 138074 800
rect 138478 0 138534 800
rect 139030 0 139086 800
rect 139490 0 139546 800
rect 139950 0 140006 800
rect 140502 0 140558 800
rect 140962 0 141018 800
rect 141422 0 141478 800
rect 141882 0 141938 800
rect 142434 0 142490 800
rect 142894 0 142950 800
rect 143354 0 143410 800
rect 143906 0 143962 800
rect 144366 0 144422 800
rect 144826 0 144882 800
rect 145378 0 145434 800
rect 145838 0 145894 800
rect 146298 0 146354 800
rect 146850 0 146906 800
rect 147310 0 147366 800
rect 147770 0 147826 800
rect 148322 0 148378 800
rect 148782 0 148838 800
rect 149242 0 149298 800
rect 149702 0 149758 800
rect 150254 0 150310 800
rect 150714 0 150770 800
rect 151174 0 151230 800
rect 151726 0 151782 800
rect 152186 0 152242 800
rect 152646 0 152702 800
rect 153198 0 153254 800
rect 153658 0 153714 800
rect 154118 0 154174 800
rect 154670 0 154726 800
rect 155130 0 155186 800
rect 155590 0 155646 800
rect 156142 0 156198 800
rect 156602 0 156658 800
rect 157062 0 157118 800
rect 157522 0 157578 800
rect 158074 0 158130 800
rect 158534 0 158590 800
rect 158994 0 159050 800
rect 159546 0 159602 800
rect 160006 0 160062 800
rect 160466 0 160522 800
rect 161018 0 161074 800
rect 161478 0 161534 800
rect 161938 0 161994 800
rect 162490 0 162546 800
rect 162950 0 163006 800
rect 163410 0 163466 800
rect 163962 0 164018 800
rect 164422 0 164478 800
rect 164882 0 164938 800
rect 165434 0 165490 800
rect 165894 0 165950 800
rect 166354 0 166410 800
rect 166814 0 166870 800
rect 167366 0 167422 800
rect 167826 0 167882 800
rect 168286 0 168342 800
rect 168838 0 168894 800
rect 169298 0 169354 800
rect 169758 0 169814 800
rect 170310 0 170366 800
rect 170770 0 170826 800
rect 171230 0 171286 800
rect 171782 0 171838 800
rect 172242 0 172298 800
rect 172702 0 172758 800
rect 173254 0 173310 800
rect 173714 0 173770 800
rect 174174 0 174230 800
rect 174634 0 174690 800
rect 175186 0 175242 800
rect 175646 0 175702 800
rect 176106 0 176162 800
rect 176658 0 176714 800
rect 177118 0 177174 800
rect 177578 0 177634 800
rect 178130 0 178186 800
rect 178590 0 178646 800
rect 179050 0 179106 800
rect 179602 0 179658 800
rect 180062 0 180118 800
rect 180522 0 180578 800
rect 181074 0 181130 800
rect 181534 0 181590 800
rect 181994 0 182050 800
rect 182454 0 182510 800
rect 183006 0 183062 800
rect 183466 0 183522 800
rect 183926 0 183982 800
rect 184478 0 184534 800
rect 184938 0 184994 800
rect 185398 0 185454 800
rect 185950 0 186006 800
rect 186410 0 186466 800
rect 186870 0 186926 800
rect 187422 0 187478 800
rect 187882 0 187938 800
rect 188342 0 188398 800
rect 188894 0 188950 800
rect 189354 0 189410 800
rect 189814 0 189870 800
rect 190366 0 190422 800
rect 190826 0 190882 800
rect 191286 0 191342 800
rect 191746 0 191802 800
rect 192298 0 192354 800
rect 192758 0 192814 800
rect 193218 0 193274 800
rect 193770 0 193826 800
rect 194230 0 194286 800
rect 194690 0 194746 800
rect 195242 0 195298 800
rect 195702 0 195758 800
rect 196162 0 196218 800
rect 196714 0 196770 800
rect 197174 0 197230 800
rect 197634 0 197690 800
rect 198186 0 198242 800
rect 198646 0 198702 800
rect 199106 0 199162 800
rect 199566 0 199622 800
rect 200118 0 200174 800
rect 200578 0 200634 800
rect 201038 0 201094 800
rect 201590 0 201646 800
rect 202050 0 202106 800
rect 202510 0 202566 800
rect 203062 0 203118 800
rect 203522 0 203578 800
rect 203982 0 204038 800
rect 204534 0 204590 800
rect 204994 0 205050 800
rect 205454 0 205510 800
rect 206006 0 206062 800
rect 206466 0 206522 800
rect 206926 0 206982 800
rect 207386 0 207442 800
rect 207938 0 207994 800
rect 208398 0 208454 800
rect 208858 0 208914 800
rect 209410 0 209466 800
rect 209870 0 209926 800
rect 210330 0 210386 800
rect 210882 0 210938 800
rect 211342 0 211398 800
rect 211802 0 211858 800
rect 212354 0 212410 800
rect 212814 0 212870 800
rect 213274 0 213330 800
rect 213826 0 213882 800
rect 214286 0 214342 800
rect 214746 0 214802 800
rect 215298 0 215354 800
rect 215758 0 215814 800
rect 216218 0 216274 800
rect 216678 0 216734 800
rect 217230 0 217286 800
rect 217690 0 217746 800
rect 218150 0 218206 800
rect 218702 0 218758 800
rect 219162 0 219218 800
rect 219622 0 219678 800
rect 220174 0 220230 800
rect 220634 0 220690 800
rect 221094 0 221150 800
rect 221646 0 221702 800
rect 222106 0 222162 800
rect 222566 0 222622 800
rect 223118 0 223174 800
rect 223578 0 223634 800
rect 224038 0 224094 800
rect 224498 0 224554 800
rect 225050 0 225106 800
rect 225510 0 225566 800
rect 225970 0 226026 800
rect 226522 0 226578 800
rect 226982 0 227038 800
rect 227442 0 227498 800
rect 227994 0 228050 800
rect 228454 0 228510 800
rect 228914 0 228970 800
rect 229466 0 229522 800
rect 229926 0 229982 800
rect 230386 0 230442 800
rect 230938 0 230994 800
rect 231398 0 231454 800
rect 231858 0 231914 800
rect 232318 0 232374 800
rect 232870 0 232926 800
rect 233330 0 233386 800
rect 233790 0 233846 800
rect 234342 0 234398 800
rect 234802 0 234858 800
rect 235262 0 235318 800
rect 235814 0 235870 800
rect 236274 0 236330 800
rect 236734 0 236790 800
rect 237286 0 237342 800
rect 237746 0 237802 800
rect 238206 0 238262 800
rect 238758 0 238814 800
rect 239218 0 239274 800
rect 239678 0 239734 800
<< obsm2 >>
rect 216 199144 974 199200
rect 1142 199144 2998 199200
rect 3166 199144 5114 199200
rect 5282 199144 7230 199200
rect 7398 199144 9254 199200
rect 9422 199144 11370 199200
rect 11538 199144 13486 199200
rect 13654 199144 15510 199200
rect 15678 199144 17626 199200
rect 17794 199144 19742 199200
rect 19910 199144 21766 199200
rect 21934 199144 23882 199200
rect 24050 199144 25998 199200
rect 26166 199144 28022 199200
rect 28190 199144 30138 199200
rect 30306 199144 32254 199200
rect 32422 199144 34278 199200
rect 34446 199144 36394 199200
rect 36562 199144 38510 199200
rect 38678 199144 40626 199200
rect 40794 199144 42650 199200
rect 42818 199144 44766 199200
rect 44934 199144 46882 199200
rect 47050 199144 48906 199200
rect 49074 199144 51022 199200
rect 51190 199144 53138 199200
rect 53306 199144 55162 199200
rect 55330 199144 57278 199200
rect 57446 199144 59394 199200
rect 59562 199144 61418 199200
rect 61586 199144 63534 199200
rect 63702 199144 65650 199200
rect 65818 199144 67674 199200
rect 67842 199144 69790 199200
rect 69958 199144 71906 199200
rect 72074 199144 74022 199200
rect 74190 199144 76046 199200
rect 76214 199144 78162 199200
rect 78330 199144 80278 199200
rect 80446 199144 82302 199200
rect 82470 199144 84418 199200
rect 84586 199144 86534 199200
rect 86702 199144 88558 199200
rect 88726 199144 90674 199200
rect 90842 199144 92790 199200
rect 92958 199144 94814 199200
rect 94982 199144 96930 199200
rect 97098 199144 99046 199200
rect 99214 199144 101070 199200
rect 101238 199144 103186 199200
rect 103354 199144 105302 199200
rect 105470 199144 107418 199200
rect 107586 199144 109442 199200
rect 109610 199144 111558 199200
rect 111726 199144 113674 199200
rect 113842 199144 115698 199200
rect 115866 199144 117814 199200
rect 117982 199144 119930 199200
rect 120098 199144 121954 199200
rect 122122 199144 124070 199200
rect 124238 199144 126186 199200
rect 126354 199144 128210 199200
rect 128378 199144 130326 199200
rect 130494 199144 132442 199200
rect 132610 199144 134466 199200
rect 134634 199144 136582 199200
rect 136750 199144 138698 199200
rect 138866 199144 140814 199200
rect 140982 199144 142838 199200
rect 143006 199144 144954 199200
rect 145122 199144 147070 199200
rect 147238 199144 149094 199200
rect 149262 199144 151210 199200
rect 151378 199144 153326 199200
rect 153494 199144 155350 199200
rect 155518 199144 157466 199200
rect 157634 199144 159582 199200
rect 159750 199144 161606 199200
rect 161774 199144 163722 199200
rect 163890 199144 165838 199200
rect 166006 199144 167862 199200
rect 168030 199144 169978 199200
rect 170146 199144 172094 199200
rect 172262 199144 174210 199200
rect 174378 199144 176234 199200
rect 176402 199144 178350 199200
rect 178518 199144 180466 199200
rect 180634 199144 182490 199200
rect 182658 199144 184606 199200
rect 184774 199144 186722 199200
rect 186890 199144 188746 199200
rect 188914 199144 190862 199200
rect 191030 199144 192978 199200
rect 193146 199144 195002 199200
rect 195170 199144 197118 199200
rect 197286 199144 199234 199200
rect 199402 199144 201258 199200
rect 201426 199144 203374 199200
rect 203542 199144 205490 199200
rect 205658 199144 207606 199200
rect 207774 199144 209630 199200
rect 209798 199144 211746 199200
rect 211914 199144 213862 199200
rect 214030 199144 215886 199200
rect 216054 199144 218002 199200
rect 218170 199144 220118 199200
rect 220286 199144 222142 199200
rect 222310 199144 224258 199200
rect 224426 199144 226374 199200
rect 226542 199144 228398 199200
rect 228566 199144 230514 199200
rect 230682 199144 232630 199200
rect 232798 199144 234654 199200
rect 234822 199144 236770 199200
rect 236938 199144 238886 199200
rect 239054 199144 239732 199200
rect 216 856 239732 199144
rect 314 2 606 856
rect 774 2 1066 856
rect 1234 2 1526 856
rect 1694 2 2078 856
rect 2246 2 2538 856
rect 2706 2 2998 856
rect 3166 2 3550 856
rect 3718 2 4010 856
rect 4178 2 4470 856
rect 4638 2 5022 856
rect 5190 2 5482 856
rect 5650 2 5942 856
rect 6110 2 6494 856
rect 6662 2 6954 856
rect 7122 2 7414 856
rect 7582 2 7966 856
rect 8134 2 8426 856
rect 8594 2 8886 856
rect 9054 2 9346 856
rect 9514 2 9898 856
rect 10066 2 10358 856
rect 10526 2 10818 856
rect 10986 2 11370 856
rect 11538 2 11830 856
rect 11998 2 12290 856
rect 12458 2 12842 856
rect 13010 2 13302 856
rect 13470 2 13762 856
rect 13930 2 14314 856
rect 14482 2 14774 856
rect 14942 2 15234 856
rect 15402 2 15786 856
rect 15954 2 16246 856
rect 16414 2 16706 856
rect 16874 2 17166 856
rect 17334 2 17718 856
rect 17886 2 18178 856
rect 18346 2 18638 856
rect 18806 2 19190 856
rect 19358 2 19650 856
rect 19818 2 20110 856
rect 20278 2 20662 856
rect 20830 2 21122 856
rect 21290 2 21582 856
rect 21750 2 22134 856
rect 22302 2 22594 856
rect 22762 2 23054 856
rect 23222 2 23606 856
rect 23774 2 24066 856
rect 24234 2 24526 856
rect 24694 2 24986 856
rect 25154 2 25538 856
rect 25706 2 25998 856
rect 26166 2 26458 856
rect 26626 2 27010 856
rect 27178 2 27470 856
rect 27638 2 27930 856
rect 28098 2 28482 856
rect 28650 2 28942 856
rect 29110 2 29402 856
rect 29570 2 29954 856
rect 30122 2 30414 856
rect 30582 2 30874 856
rect 31042 2 31426 856
rect 31594 2 31886 856
rect 32054 2 32346 856
rect 32514 2 32898 856
rect 33066 2 33358 856
rect 33526 2 33818 856
rect 33986 2 34278 856
rect 34446 2 34830 856
rect 34998 2 35290 856
rect 35458 2 35750 856
rect 35918 2 36302 856
rect 36470 2 36762 856
rect 36930 2 37222 856
rect 37390 2 37774 856
rect 37942 2 38234 856
rect 38402 2 38694 856
rect 38862 2 39246 856
rect 39414 2 39706 856
rect 39874 2 40166 856
rect 40334 2 40718 856
rect 40886 2 41178 856
rect 41346 2 41638 856
rect 41806 2 42098 856
rect 42266 2 42650 856
rect 42818 2 43110 856
rect 43278 2 43570 856
rect 43738 2 44122 856
rect 44290 2 44582 856
rect 44750 2 45042 856
rect 45210 2 45594 856
rect 45762 2 46054 856
rect 46222 2 46514 856
rect 46682 2 47066 856
rect 47234 2 47526 856
rect 47694 2 47986 856
rect 48154 2 48538 856
rect 48706 2 48998 856
rect 49166 2 49458 856
rect 49626 2 49918 856
rect 50086 2 50470 856
rect 50638 2 50930 856
rect 51098 2 51390 856
rect 51558 2 51942 856
rect 52110 2 52402 856
rect 52570 2 52862 856
rect 53030 2 53414 856
rect 53582 2 53874 856
rect 54042 2 54334 856
rect 54502 2 54886 856
rect 55054 2 55346 856
rect 55514 2 55806 856
rect 55974 2 56358 856
rect 56526 2 56818 856
rect 56986 2 57278 856
rect 57446 2 57830 856
rect 57998 2 58290 856
rect 58458 2 58750 856
rect 58918 2 59210 856
rect 59378 2 59762 856
rect 59930 2 60222 856
rect 60390 2 60682 856
rect 60850 2 61234 856
rect 61402 2 61694 856
rect 61862 2 62154 856
rect 62322 2 62706 856
rect 62874 2 63166 856
rect 63334 2 63626 856
rect 63794 2 64178 856
rect 64346 2 64638 856
rect 64806 2 65098 856
rect 65266 2 65650 856
rect 65818 2 66110 856
rect 66278 2 66570 856
rect 66738 2 67030 856
rect 67198 2 67582 856
rect 67750 2 68042 856
rect 68210 2 68502 856
rect 68670 2 69054 856
rect 69222 2 69514 856
rect 69682 2 69974 856
rect 70142 2 70526 856
rect 70694 2 70986 856
rect 71154 2 71446 856
rect 71614 2 71998 856
rect 72166 2 72458 856
rect 72626 2 72918 856
rect 73086 2 73470 856
rect 73638 2 73930 856
rect 74098 2 74390 856
rect 74558 2 74850 856
rect 75018 2 75402 856
rect 75570 2 75862 856
rect 76030 2 76322 856
rect 76490 2 76874 856
rect 77042 2 77334 856
rect 77502 2 77794 856
rect 77962 2 78346 856
rect 78514 2 78806 856
rect 78974 2 79266 856
rect 79434 2 79818 856
rect 79986 2 80278 856
rect 80446 2 80738 856
rect 80906 2 81290 856
rect 81458 2 81750 856
rect 81918 2 82210 856
rect 82378 2 82762 856
rect 82930 2 83222 856
rect 83390 2 83682 856
rect 83850 2 84142 856
rect 84310 2 84694 856
rect 84862 2 85154 856
rect 85322 2 85614 856
rect 85782 2 86166 856
rect 86334 2 86626 856
rect 86794 2 87086 856
rect 87254 2 87638 856
rect 87806 2 88098 856
rect 88266 2 88558 856
rect 88726 2 89110 856
rect 89278 2 89570 856
rect 89738 2 90030 856
rect 90198 2 90582 856
rect 90750 2 91042 856
rect 91210 2 91502 856
rect 91670 2 91962 856
rect 92130 2 92514 856
rect 92682 2 92974 856
rect 93142 2 93434 856
rect 93602 2 93986 856
rect 94154 2 94446 856
rect 94614 2 94906 856
rect 95074 2 95458 856
rect 95626 2 95918 856
rect 96086 2 96378 856
rect 96546 2 96930 856
rect 97098 2 97390 856
rect 97558 2 97850 856
rect 98018 2 98402 856
rect 98570 2 98862 856
rect 99030 2 99322 856
rect 99490 2 99782 856
rect 99950 2 100334 856
rect 100502 2 100794 856
rect 100962 2 101254 856
rect 101422 2 101806 856
rect 101974 2 102266 856
rect 102434 2 102726 856
rect 102894 2 103278 856
rect 103446 2 103738 856
rect 103906 2 104198 856
rect 104366 2 104750 856
rect 104918 2 105210 856
rect 105378 2 105670 856
rect 105838 2 106222 856
rect 106390 2 106682 856
rect 106850 2 107142 856
rect 107310 2 107694 856
rect 107862 2 108154 856
rect 108322 2 108614 856
rect 108782 2 109074 856
rect 109242 2 109626 856
rect 109794 2 110086 856
rect 110254 2 110546 856
rect 110714 2 111098 856
rect 111266 2 111558 856
rect 111726 2 112018 856
rect 112186 2 112570 856
rect 112738 2 113030 856
rect 113198 2 113490 856
rect 113658 2 114042 856
rect 114210 2 114502 856
rect 114670 2 114962 856
rect 115130 2 115514 856
rect 115682 2 115974 856
rect 116142 2 116434 856
rect 116602 2 116894 856
rect 117062 2 117446 856
rect 117614 2 117906 856
rect 118074 2 118366 856
rect 118534 2 118918 856
rect 119086 2 119378 856
rect 119546 2 119838 856
rect 120006 2 120390 856
rect 120558 2 120850 856
rect 121018 2 121310 856
rect 121478 2 121862 856
rect 122030 2 122322 856
rect 122490 2 122782 856
rect 122950 2 123334 856
rect 123502 2 123794 856
rect 123962 2 124254 856
rect 124422 2 124714 856
rect 124882 2 125266 856
rect 125434 2 125726 856
rect 125894 2 126186 856
rect 126354 2 126738 856
rect 126906 2 127198 856
rect 127366 2 127658 856
rect 127826 2 128210 856
rect 128378 2 128670 856
rect 128838 2 129130 856
rect 129298 2 129682 856
rect 129850 2 130142 856
rect 130310 2 130602 856
rect 130770 2 131154 856
rect 131322 2 131614 856
rect 131782 2 132074 856
rect 132242 2 132534 856
rect 132702 2 133086 856
rect 133254 2 133546 856
rect 133714 2 134006 856
rect 134174 2 134558 856
rect 134726 2 135018 856
rect 135186 2 135478 856
rect 135646 2 136030 856
rect 136198 2 136490 856
rect 136658 2 136950 856
rect 137118 2 137502 856
rect 137670 2 137962 856
rect 138130 2 138422 856
rect 138590 2 138974 856
rect 139142 2 139434 856
rect 139602 2 139894 856
rect 140062 2 140446 856
rect 140614 2 140906 856
rect 141074 2 141366 856
rect 141534 2 141826 856
rect 141994 2 142378 856
rect 142546 2 142838 856
rect 143006 2 143298 856
rect 143466 2 143850 856
rect 144018 2 144310 856
rect 144478 2 144770 856
rect 144938 2 145322 856
rect 145490 2 145782 856
rect 145950 2 146242 856
rect 146410 2 146794 856
rect 146962 2 147254 856
rect 147422 2 147714 856
rect 147882 2 148266 856
rect 148434 2 148726 856
rect 148894 2 149186 856
rect 149354 2 149646 856
rect 149814 2 150198 856
rect 150366 2 150658 856
rect 150826 2 151118 856
rect 151286 2 151670 856
rect 151838 2 152130 856
rect 152298 2 152590 856
rect 152758 2 153142 856
rect 153310 2 153602 856
rect 153770 2 154062 856
rect 154230 2 154614 856
rect 154782 2 155074 856
rect 155242 2 155534 856
rect 155702 2 156086 856
rect 156254 2 156546 856
rect 156714 2 157006 856
rect 157174 2 157466 856
rect 157634 2 158018 856
rect 158186 2 158478 856
rect 158646 2 158938 856
rect 159106 2 159490 856
rect 159658 2 159950 856
rect 160118 2 160410 856
rect 160578 2 160962 856
rect 161130 2 161422 856
rect 161590 2 161882 856
rect 162050 2 162434 856
rect 162602 2 162894 856
rect 163062 2 163354 856
rect 163522 2 163906 856
rect 164074 2 164366 856
rect 164534 2 164826 856
rect 164994 2 165378 856
rect 165546 2 165838 856
rect 166006 2 166298 856
rect 166466 2 166758 856
rect 166926 2 167310 856
rect 167478 2 167770 856
rect 167938 2 168230 856
rect 168398 2 168782 856
rect 168950 2 169242 856
rect 169410 2 169702 856
rect 169870 2 170254 856
rect 170422 2 170714 856
rect 170882 2 171174 856
rect 171342 2 171726 856
rect 171894 2 172186 856
rect 172354 2 172646 856
rect 172814 2 173198 856
rect 173366 2 173658 856
rect 173826 2 174118 856
rect 174286 2 174578 856
rect 174746 2 175130 856
rect 175298 2 175590 856
rect 175758 2 176050 856
rect 176218 2 176602 856
rect 176770 2 177062 856
rect 177230 2 177522 856
rect 177690 2 178074 856
rect 178242 2 178534 856
rect 178702 2 178994 856
rect 179162 2 179546 856
rect 179714 2 180006 856
rect 180174 2 180466 856
rect 180634 2 181018 856
rect 181186 2 181478 856
rect 181646 2 181938 856
rect 182106 2 182398 856
rect 182566 2 182950 856
rect 183118 2 183410 856
rect 183578 2 183870 856
rect 184038 2 184422 856
rect 184590 2 184882 856
rect 185050 2 185342 856
rect 185510 2 185894 856
rect 186062 2 186354 856
rect 186522 2 186814 856
rect 186982 2 187366 856
rect 187534 2 187826 856
rect 187994 2 188286 856
rect 188454 2 188838 856
rect 189006 2 189298 856
rect 189466 2 189758 856
rect 189926 2 190310 856
rect 190478 2 190770 856
rect 190938 2 191230 856
rect 191398 2 191690 856
rect 191858 2 192242 856
rect 192410 2 192702 856
rect 192870 2 193162 856
rect 193330 2 193714 856
rect 193882 2 194174 856
rect 194342 2 194634 856
rect 194802 2 195186 856
rect 195354 2 195646 856
rect 195814 2 196106 856
rect 196274 2 196658 856
rect 196826 2 197118 856
rect 197286 2 197578 856
rect 197746 2 198130 856
rect 198298 2 198590 856
rect 198758 2 199050 856
rect 199218 2 199510 856
rect 199678 2 200062 856
rect 200230 2 200522 856
rect 200690 2 200982 856
rect 201150 2 201534 856
rect 201702 2 201994 856
rect 202162 2 202454 856
rect 202622 2 203006 856
rect 203174 2 203466 856
rect 203634 2 203926 856
rect 204094 2 204478 856
rect 204646 2 204938 856
rect 205106 2 205398 856
rect 205566 2 205950 856
rect 206118 2 206410 856
rect 206578 2 206870 856
rect 207038 2 207330 856
rect 207498 2 207882 856
rect 208050 2 208342 856
rect 208510 2 208802 856
rect 208970 2 209354 856
rect 209522 2 209814 856
rect 209982 2 210274 856
rect 210442 2 210826 856
rect 210994 2 211286 856
rect 211454 2 211746 856
rect 211914 2 212298 856
rect 212466 2 212758 856
rect 212926 2 213218 856
rect 213386 2 213770 856
rect 213938 2 214230 856
rect 214398 2 214690 856
rect 214858 2 215242 856
rect 215410 2 215702 856
rect 215870 2 216162 856
rect 216330 2 216622 856
rect 216790 2 217174 856
rect 217342 2 217634 856
rect 217802 2 218094 856
rect 218262 2 218646 856
rect 218814 2 219106 856
rect 219274 2 219566 856
rect 219734 2 220118 856
rect 220286 2 220578 856
rect 220746 2 221038 856
rect 221206 2 221590 856
rect 221758 2 222050 856
rect 222218 2 222510 856
rect 222678 2 223062 856
rect 223230 2 223522 856
rect 223690 2 223982 856
rect 224150 2 224442 856
rect 224610 2 224994 856
rect 225162 2 225454 856
rect 225622 2 225914 856
rect 226082 2 226466 856
rect 226634 2 226926 856
rect 227094 2 227386 856
rect 227554 2 227938 856
rect 228106 2 228398 856
rect 228566 2 228858 856
rect 229026 2 229410 856
rect 229578 2 229870 856
rect 230038 2 230330 856
rect 230498 2 230882 856
rect 231050 2 231342 856
rect 231510 2 231802 856
rect 231970 2 232262 856
rect 232430 2 232814 856
rect 232982 2 233274 856
rect 233442 2 233734 856
rect 233902 2 234286 856
rect 234454 2 234746 856
rect 234914 2 235206 856
rect 235374 2 235758 856
rect 235926 2 236218 856
rect 236386 2 236678 856
rect 236846 2 237230 856
rect 237398 2 237690 856
rect 237858 2 238150 856
rect 238318 2 238702 856
rect 238870 2 239162 856
rect 239330 2 239622 856
<< metal3 >>
rect 0 99968 800 100088
<< obsm3 >>
rect 800 100168 237899 197505
rect 880 99888 237899 100168
rect 800 35 237899 99888
<< metal4 >>
rect 4208 2128 4528 197520
rect 4868 2176 5188 197472
rect 5528 2176 5848 197472
rect 6188 2176 6508 197472
rect 19568 2128 19888 197520
rect 20228 2176 20548 197472
rect 20888 2176 21208 197472
rect 21548 2176 21868 197472
rect 34928 2128 35248 197520
rect 35588 2176 35908 197472
rect 36248 2176 36568 197472
rect 36908 2176 37228 197472
rect 50288 2128 50608 197520
rect 50948 2176 51268 197472
rect 51608 2176 51928 197472
rect 52268 2176 52588 197472
rect 65648 2128 65968 197520
rect 66308 2176 66628 197472
rect 66968 2176 67288 197472
rect 67628 2176 67948 197472
rect 81008 2128 81328 197520
rect 81668 2176 81988 197472
rect 82328 2176 82648 197472
rect 82988 2176 83308 197472
rect 96368 2128 96688 197520
rect 97028 2176 97348 197472
rect 97688 2176 98008 197472
rect 98348 2176 98668 197472
rect 111728 2128 112048 197520
rect 112388 2176 112708 197472
rect 113048 2176 113368 197472
rect 113708 2176 114028 197472
rect 127088 2128 127408 197520
rect 127748 2176 128068 197472
rect 128408 2176 128728 197472
rect 129068 2176 129388 197472
rect 142448 2128 142768 197520
rect 143108 2176 143428 197472
rect 143768 2176 144088 197472
rect 144428 2176 144748 197472
rect 157808 2128 158128 197520
rect 158468 2176 158788 197472
rect 159128 2176 159448 197472
rect 159788 2176 160108 197472
rect 173168 2128 173488 197520
rect 173828 2176 174148 197472
rect 174488 2176 174808 197472
rect 175148 2176 175468 197472
rect 188528 2128 188848 197520
rect 189188 2176 189508 197472
rect 189848 2176 190168 197472
rect 190508 2176 190828 197472
rect 203888 2128 204208 197520
rect 204548 2176 204868 197472
rect 205208 2176 205528 197472
rect 205868 2176 206188 197472
rect 219248 2128 219568 197520
rect 219908 2176 220228 197472
rect 220568 2176 220888 197472
rect 221228 2176 221548 197472
rect 234608 2128 234928 197520
rect 235268 2176 235588 197472
rect 235928 2176 236248 197472
rect 236588 2176 236908 197472
<< obsm4 >>
rect 124627 2048 127008 22269
rect 127488 2096 127668 22269
rect 128148 2096 128328 22269
rect 128808 2096 128988 22269
rect 129468 2096 142368 22269
rect 127488 2048 142368 2096
rect 142848 2096 143028 22269
rect 143508 2096 143688 22269
rect 144168 2096 144348 22269
rect 144828 2096 157728 22269
rect 142848 2048 157728 2096
rect 158208 2096 158388 22269
rect 158868 2096 159048 22269
rect 159528 2096 159708 22269
rect 160188 2096 173088 22269
rect 158208 2048 173088 2096
rect 173568 2096 173748 22269
rect 174228 2096 174408 22269
rect 174888 2096 175068 22269
rect 175548 2096 188448 22269
rect 173568 2048 188448 2096
rect 188928 2096 189108 22269
rect 189588 2096 189768 22269
rect 190248 2096 190428 22269
rect 190908 2096 195901 22269
rect 188928 2048 195901 2096
rect 124627 443 195901 2048
<< labels >>
rlabel metal2 s 1030 199200 1086 200000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 63590 199200 63646 200000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 69846 199200 69902 200000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 76102 199200 76158 200000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 82358 199200 82414 200000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 88614 199200 88670 200000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 94870 199200 94926 200000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 101126 199200 101182 200000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 107474 199200 107530 200000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 113730 199200 113786 200000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 119986 199200 120042 200000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7286 199200 7342 200000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 126242 199200 126298 200000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 132498 199200 132554 200000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 138754 199200 138810 200000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 145010 199200 145066 200000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 151266 199200 151322 200000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 157522 199200 157578 200000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 163778 199200 163834 200000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 170034 199200 170090 200000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 176290 199200 176346 200000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 182546 199200 182602 200000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 13542 199200 13598 200000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 188802 199200 188858 200000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 195058 199200 195114 200000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 201314 199200 201370 200000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 207662 199200 207718 200000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 213918 199200 213974 200000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 220174 199200 220230 200000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 226430 199200 226486 200000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 232686 199200 232742 200000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 19798 199200 19854 200000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 26054 199200 26110 200000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 32310 199200 32366 200000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 38566 199200 38622 200000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 44822 199200 44878 200000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 51078 199200 51134 200000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 57334 199200 57390 200000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3054 199200 3110 200000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 65706 199200 65762 200000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 71962 199200 72018 200000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 78218 199200 78274 200000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 84474 199200 84530 200000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 90730 199200 90786 200000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 96986 199200 97042 200000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 103242 199200 103298 200000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 109498 199200 109554 200000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 115754 199200 115810 200000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 122010 199200 122066 200000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9310 199200 9366 200000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 128266 199200 128322 200000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 134522 199200 134578 200000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 140870 199200 140926 200000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 147126 199200 147182 200000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 153382 199200 153438 200000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 159638 199200 159694 200000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 165894 199200 165950 200000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 172150 199200 172206 200000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 178406 199200 178462 200000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 184662 199200 184718 200000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 15566 199200 15622 200000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 190918 199200 190974 200000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 197174 199200 197230 200000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 203430 199200 203486 200000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 209686 199200 209742 200000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 215942 199200 215998 200000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 222198 199200 222254 200000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 228454 199200 228510 200000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 234710 199200 234766 200000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 21822 199200 21878 200000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 28078 199200 28134 200000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 34334 199200 34390 200000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 40682 199200 40738 200000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 46938 199200 46994 200000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 53194 199200 53250 200000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 59450 199200 59506 200000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 5170 199200 5226 200000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 67730 199200 67786 200000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 74078 199200 74134 200000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 80334 199200 80390 200000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 86590 199200 86646 200000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 92846 199200 92902 200000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 99102 199200 99158 200000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 105358 199200 105414 200000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 111614 199200 111670 200000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 117870 199200 117926 200000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 124126 199200 124182 200000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11426 199200 11482 200000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 130382 199200 130438 200000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 136638 199200 136694 200000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 142894 199200 142950 200000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 149150 199200 149206 200000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 155406 199200 155462 200000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 161662 199200 161718 200000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 167918 199200 167974 200000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 174266 199200 174322 200000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 180522 199200 180578 200000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 186778 199200 186834 200000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 17682 199200 17738 200000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 193034 199200 193090 200000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 199290 199200 199346 200000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 205546 199200 205602 200000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 211802 199200 211858 200000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 218058 199200 218114 200000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 224314 199200 224370 200000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 230570 199200 230626 200000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 236826 199200 236882 200000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 23938 199200 23994 200000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 30194 199200 30250 200000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 36450 199200 36506 200000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 42706 199200 42762 200000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 48962 199200 49018 200000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 55218 199200 55274 200000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 61474 199200 61530 200000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 239678 0 239734 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 238942 199200 238998 200000 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 51998 0 52054 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 198646 0 198702 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 200118 0 200174 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 203062 0 203118 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 204534 0 204590 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 206006 0 206062 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 207386 0 207442 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 208858 0 208914 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 210330 0 210386 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 213274 0 213330 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 216218 0 216274 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 217690 0 217746 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 219162 0 219218 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 220634 0 220690 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 222106 0 222162 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 223578 0 223634 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 226522 0 226578 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 227994 0 228050 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 229466 0 229522 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 230938 0 230994 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 232318 0 232374 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 233790 0 233846 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 235262 0 235318 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 236734 0 236790 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 238206 0 238262 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 73986 0 74042 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 87142 0 87198 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 90086 0 90142 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 104806 0 104862 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 116490 0 116546 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 119434 0 119490 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 122378 0 122434 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 128266 0 128322 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 132590 0 132646 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 142894 0 142950 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 144366 0 144422 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 161938 0 161994 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 167826 0 167882 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 173714 0 173770 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 175186 0 175242 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 179602 0 179658 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 181074 0 181130 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 182454 0 182510 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 183926 0 183982 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 185398 0 185454 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 186870 0 186926 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 189814 0 189870 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 191286 0 191342 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 192758 0 192814 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 194230 0 194286 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 195702 0 195758 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 197174 0 197230 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 199106 0 199162 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 202050 0 202106 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 203522 0 203578 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 204994 0 205050 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 206466 0 206522 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 207938 0 207994 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 209410 0 209466 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 210882 0 210938 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 212354 0 212410 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 213826 0 213882 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 215298 0 215354 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 216678 0 216734 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 218150 0 218206 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 219622 0 219678 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 221094 0 221150 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 222566 0 222622 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 224038 0 224094 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 225510 0 225566 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 226982 0 227038 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 68558 0 68614 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 228454 0 228510 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 229926 0 229982 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 231398 0 231454 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 232870 0 232926 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 234342 0 234398 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 235814 0 235870 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 237286 0 237342 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 238758 0 238814 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 70030 0 70086 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 72974 0 73030 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 74446 0 74502 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 77390 0 77446 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 80334 0 80390 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 81806 0 81862 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 83278 0 83334 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 84750 0 84806 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 87694 0 87750 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 92018 0 92074 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 93490 0 93546 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 94962 0 95018 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 55402 0 55458 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 97906 0 97962 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 102322 0 102378 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 111154 0 111210 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 116950 0 117006 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 127254 0 127310 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 128726 0 128782 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 140502 0 140558 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 143354 0 143410 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 144826 0 144882 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 61290 0 61346 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 155130 0 155186 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 156602 0 156658 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 165434 0 165490 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 168286 0 168342 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 171230 0 171286 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 172702 0 172758 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 175646 0 175702 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 177118 0 177174 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 178590 0 178646 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 180062 0 180118 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 181534 0 181590 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 183006 0 183062 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 64234 0 64290 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 184478 0 184534 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 185950 0 186006 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 187422 0 187478 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 188894 0 188950 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 190366 0 190422 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 191746 0 191802 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 194690 0 194746 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 196162 0 196218 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 197634 0 197690 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 65706 0 65762 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 199566 0 199622 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 201038 0 201094 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 202510 0 202566 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 203982 0 204038 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 205454 0 205510 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 206926 0 206982 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 209870 0 209926 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 211342 0 211398 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 214286 0 214342 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 215758 0 215814 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 217230 0 217286 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 218702 0 218758 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 220174 0 220230 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 221646 0 221702 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 224498 0 224554 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 225970 0 226026 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 227442 0 227498 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 230386 0 230442 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 231858 0 231914 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 233330 0 233386 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 234802 0 234858 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 236274 0 236330 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 237746 0 237802 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 239218 0 239274 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 74906 0 74962 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 54390 0 54446 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 83738 0 83794 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 98458 0 98514 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 120446 0 120502 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 145378 0 145434 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 154118 0 154174 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 158534 0 158590 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 161478 0 161534 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 164422 0 164478 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 173254 0 173310 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 174634 0 174690 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 177578 0 177634 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 179050 0 179106 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 181994 0 182050 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 184938 0 184994 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 189354 0 189410 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 190826 0 190882 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 192298 0 192354 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 193770 0 193826 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 195242 0 195298 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 196714 0 196770 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 202 0 258 800 6 wb_clk_i
port 502 nsew signal input
rlabel metal2 s 662 0 718 800 6 wb_rst_i
port 503 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 wbs_ack_o
port 504 nsew signal output
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[0]
port 505 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[10]
port 506 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_adr_i[11]
port 507 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[12]
port 508 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[13]
port 509 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_adr_i[14]
port 510 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 wbs_adr_i[15]
port 511 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_adr_i[16]
port 512 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[17]
port 513 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 wbs_adr_i[18]
port 514 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[19]
port 515 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_adr_i[1]
port 516 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wbs_adr_i[20]
port 517 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[21]
port 518 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 wbs_adr_i[22]
port 519 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_adr_i[23]
port 520 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_adr_i[24]
port 521 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_adr_i[25]
port 522 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[26]
port 523 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[27]
port 524 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 wbs_adr_i[28]
port 525 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[29]
port 526 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_adr_i[2]
port 527 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 wbs_adr_i[30]
port 528 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[31]
port 529 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_adr_i[3]
port 530 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[4]
port 531 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[5]
port 532 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[6]
port 533 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_adr_i[7]
port 534 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_adr_i[8]
port 535 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[9]
port 536 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_cyc_i
port 537 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_i[0]
port 538 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_i[10]
port 539 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[11]
port 540 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[12]
port 541 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_i[13]
port 542 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[14]
port 543 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[15]
port 544 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[16]
port 545 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[17]
port 546 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[18]
port 547 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_dat_i[19]
port 548 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_i[1]
port 549 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[20]
port 550 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[21]
port 551 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[22]
port 552 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_i[23]
port 553 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_i[24]
port 554 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[25]
port 555 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[26]
port 556 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_i[27]
port 557 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[28]
port 558 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[29]
port 559 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[2]
port 560 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_i[30]
port 561 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_i[31]
port 562 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[3]
port 563 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[4]
port 564 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[5]
port 565 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_i[6]
port 566 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[7]
port 567 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_dat_i[8]
port 568 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[9]
port 569 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_dat_o[0]
port 570 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[10]
port 571 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_o[11]
port 572 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[12]
port 573 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 wbs_dat_o[13]
port 574 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_o[14]
port 575 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[15]
port 576 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_o[16]
port 577 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 wbs_dat_o[17]
port 578 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 wbs_dat_o[18]
port 579 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_o[19]
port 580 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[1]
port 581 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 wbs_dat_o[20]
port 582 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[21]
port 583 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_o[22]
port 584 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 wbs_dat_o[23]
port 585 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 wbs_dat_o[24]
port 586 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[25]
port 587 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[26]
port 588 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[27]
port 589 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_o[28]
port 590 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[29]
port 591 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_dat_o[2]
port 592 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_o[30]
port 593 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_o[31]
port 594 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[3]
port 595 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[4]
port 596 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[5]
port 597 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_o[6]
port 598 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[7]
port 599 nsew signal output
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_o[8]
port 600 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[9]
port 601 nsew signal output
rlabel metal2 s 4526 0 4582 800 6 wbs_sel_i[0]
port 602 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_sel_i[1]
port 603 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_sel_i[2]
port 604 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 wbs_sel_i[3]
port 605 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_stb_i
port 606 nsew signal input
rlabel metal2 s 2594 0 2650 800 6 wbs_we_i
port 607 nsew signal input
rlabel metal4 s 219248 2128 219568 197520 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 609 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 610 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 611 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 612 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 613 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 614 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 615 nsew power bidirectional
rlabel metal4 s 234608 2128 234928 197520 6 vssd1
port 616 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 197520 6 vssd1
port 617 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 618 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 619 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 620 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 621 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 622 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 623 nsew ground bidirectional
rlabel metal4 s 219908 2176 220228 197472 6 vccd2
port 624 nsew power bidirectional
rlabel metal4 s 189188 2176 189508 197472 6 vccd2
port 625 nsew power bidirectional
rlabel metal4 s 158468 2176 158788 197472 6 vccd2
port 626 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 197472 6 vccd2
port 627 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 197472 6 vccd2
port 628 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 197472 6 vccd2
port 629 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 197472 6 vccd2
port 630 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 197472 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 235268 2176 235588 197472 6 vssd2
port 632 nsew ground bidirectional
rlabel metal4 s 204548 2176 204868 197472 6 vssd2
port 633 nsew ground bidirectional
rlabel metal4 s 173828 2176 174148 197472 6 vssd2
port 634 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 197472 6 vssd2
port 635 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 197472 6 vssd2
port 636 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 197472 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 197472 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 197472 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 220568 2176 220888 197472 6 vdda1
port 640 nsew power bidirectional
rlabel metal4 s 189848 2176 190168 197472 6 vdda1
port 641 nsew power bidirectional
rlabel metal4 s 159128 2176 159448 197472 6 vdda1
port 642 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 197472 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 197472 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 197472 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 197472 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 197472 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 235928 2176 236248 197472 6 vssa1
port 648 nsew ground bidirectional
rlabel metal4 s 205208 2176 205528 197472 6 vssa1
port 649 nsew ground bidirectional
rlabel metal4 s 174488 2176 174808 197472 6 vssa1
port 650 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 197472 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 197472 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 197472 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 197472 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 197472 6 vssa1
port 655 nsew ground bidirectional
rlabel metal4 s 221228 2176 221548 197472 6 vdda2
port 656 nsew power bidirectional
rlabel metal4 s 190508 2176 190828 197472 6 vdda2
port 657 nsew power bidirectional
rlabel metal4 s 159788 2176 160108 197472 6 vdda2
port 658 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 197472 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 197472 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 197472 6 vdda2
port 661 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 197472 6 vdda2
port 662 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 197472 6 vdda2
port 663 nsew power bidirectional
rlabel metal4 s 236588 2176 236908 197472 6 vssa2
port 664 nsew ground bidirectional
rlabel metal4 s 205868 2176 206188 197472 6 vssa2
port 665 nsew ground bidirectional
rlabel metal4 s 175148 2176 175468 197472 6 vssa2
port 666 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 197472 6 vssa2
port 667 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 197472 6 vssa2
port 668 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 197472 6 vssa2
port 669 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 197472 6 vssa2
port 670 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 197472 6 vssa2
port 671 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 240000 200000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj_example/runs/user_proj_example/results/magic/user_proj_example.gds
string GDS_END 32758296
string GDS_START 601002
<< end >>

